`default_nettype none

module pipe_fwd_controller(
    input EXE_wreg,
    input EXE_m2reg, 
    input [4: 0] ID_rs, 
    input [4: 0] ID_rt, 
    input [4: 0] EXE_write_reg_number, 

    
);
    // 直通处理器

    

endmodule